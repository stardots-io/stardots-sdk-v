module stardots

// SDK version
pub const sdk_version = '1.0.0'

// Endpoint Request the endpoint of the stardots server.
pub const endpoint = 'https://api.stardots.io'

// Default request timeout, unit: seconds
pub const default_request_timeout = 30 